module sevenseg2seven(ledsegments,hex0,hex1,hex2,hex3,hex4,hex5,hex6);
	input [3:0] data;
	output ledsegments;
	reg [6:0] ledsegments;
endmodule